module not_1in_v (
  input A,
  output Z
  );

  not(Z, A);

endmodule // not_1in_v
