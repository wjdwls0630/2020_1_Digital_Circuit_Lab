module bit8_adder_tb ();
  reg Cin;
  reg [7:0] A;
  reg [7:0] B;
  initial begin
    Cin <= 1'b0;
    A <= 8'b0;
    B <= 8'b0;
  end

  initial begin
    #10 A <= 8'b01010101;
    B <= 8'b01010101;
    #10 A <= 8'b01010101;
    B <= 8'b10101010;
    #10 A <= 8'b10101010;
    B <= 8'b10101010;
    #10 A <= 8'b00110011;
    B <= 8'b00110011;
    #10 A <= 8'b00110011;
    B <= 8'b11001100;
    #10 A <= 8'b11001100;
    B <= 8'b11001100;
    #10 A <= 8'b00001111;
    B <= 8'b00001111;
    #10 A <= 8'b00001111;
    B <= 8'b11110000;
    #10 A <= 8'b11110000;
    B <= 8'b11110000;
    #10 A <= 8'b00000000;
    B <= 8'b00001111;
    #10 A <= 8'b11111111; //12
    B <= 8'b00000000;
    #10 A <= 8'b01111111; //13
    B <= 8'b11111111;
    #10 A <= 8'b11111111;
    B <= 8'b11111111; // 14

    #10 A <= 8'b00000000;
    B <= 8'b00000000;
    Cin <= 1'b1;
    #10 A <= 8'b01010101;
    B <= 8'b01010101;
    #10 A <= 8'b01010101;
    B <= 8'b10101010;
    #10 A <= 8'b10101010;
    B <= 8'b10101010;
    #10 A <= 8'b00110011;
    B <= 8'b00110011;
    #10 A <= 8'b00110011;
    B <= 8'b11001100;
    #10 A <= 8'b11001100;
    B <= 8'b11001100;
    #10 A <= 8'b00001111;
    B <= 8'b00001111;
    #10 A <= 8'b00001111;
    B <= 8'b11110000;
    #10 A <= 8'b11110000;
    B <= 8'b11110000;
    #10 A <= 8'b00000000;
    B <= 8'b00001111;
    #10 A <= 8'b11111111; //12
    B <= 8'b00000000;
    #10 A <= 8'b01111111; //13
    B <= 8'b11111111;
    #10 A <= 8'b11111111;
    B <= 8'b11111111; // 14
  end
  wire [7:0] S;
  wire Cout;
  always @ ( S, Cout ) begin
    $monitor("%8b %b", S, Cout);
  end
  bit8_adder_v bit8_adder_v(
    .A(A),
    .B(B),
    .Cin(Cin),
    .S(S),
    .Cout(Cout)
  );


endmodule //multiplexer_8to1_tb
